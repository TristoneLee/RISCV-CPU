module FetchBuffer(input wire clk,
                   input wire [31:0] _PC,
                   output wire [31:0] d_out);
    
    
    
    
endmodule
